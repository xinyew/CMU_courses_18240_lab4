`default_nettype none

module bus_memory();
    bus
    memory
endmodule: memory